`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2017/12/30 13:38:08
// Design Name: 
// Module Name: VGA_char
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module VGA_char(
    input [2:0] dH,
    input [3:0] dV,
    input [5:0] alph,
    input [9:0] dcnt,
    output reg Point
    );
    reg [127:0] Char_Matrix[53:0];
    initial
    begin
        Char_Matrix[0] = {8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00}; // space
        Char_Matrix[1] = {8'h00,8'h00,8'h08,8'h1C,8'h36,8'h63,8'h63,8'h63,8'h7F,8'h63,8'h63,8'h63,8'h00,8'h00,8'h00,8'h00}; // A
        Char_Matrix[2] = {8'h00,8'h00,8'h7E,8'h33,8'h33,8'h33,8'h3E,8'h33,8'h33,8'h33,8'h33,8'h7E,8'h00,8'h00,8'h00,8'h00}; // B
        Char_Matrix[3] = {8'h00,8'h00,8'h1E,8'h33,8'h61,8'h60,8'h60,8'h60,8'h60,8'h61,8'h33,8'h1E,8'h00,8'h00,8'h00,8'h00}; // C
        Char_Matrix[4] = {8'h00,8'h00,8'h7C,8'h36,8'h33,8'h33,8'h33,8'h33,8'h33,8'h33,8'h36,8'h7C,8'h00,8'h00,8'h00,8'h00}; // D
        Char_Matrix[5] = {8'h00,8'h00,8'h7F,8'h33,8'h31,8'h34,8'h3C,8'h34,8'h30,8'h31,8'h33,8'h7F,8'h00,8'h00,8'h00,8'h00}; // E
        Char_Matrix[6] = {8'h00,8'h00,8'h7F,8'h33,8'h31,8'h34,8'h3C,8'h34,8'h30,8'h30,8'h30,8'h78,8'h00,8'h00,8'h00,8'h00}; // F
        Char_Matrix[7] = {8'h00,8'h00,8'h1E,8'h33,8'h61,8'h60,8'h60,8'h6F,8'h63,8'h63,8'h37,8'h1D,8'h00,8'h00,8'h00,8'h00}; // G
        Char_Matrix[8] = {8'h00,8'h00,8'h63,8'h63,8'h63,8'h63,8'h7F,8'h63,8'h63,8'h63,8'h63,8'h63,8'h00,8'h00,8'h00,8'h00}; // H
        Char_Matrix[9] = {8'h00,8'h00,8'h3C,8'h18,8'h18,8'h18,8'h18,8'h18,8'h18,8'h18,8'h18,8'h3C,8'h00,8'h00,8'h00,8'h00}; // I
        Char_Matrix[10] = {8'h00,8'h00,8'h0F,8'h06,8'h06,8'h06,8'h06,8'h06,8'h06,8'h66,8'h66,8'h3C,8'h00,8'h00,8'h00,8'h00}; // J
        Char_Matrix[11] = {8'h00,8'h00,8'h73,8'h33,8'h36,8'h36,8'h3C,8'h36,8'h36,8'h33,8'h33,8'h73,8'h00,8'h00,8'h00,8'h00}; // K
        Char_Matrix[12] = {8'h00,8'h00,8'h78,8'h30,8'h30,8'h30,8'h30,8'h30,8'h30,8'h31,8'h33,8'h7F,8'h00,8'h00,8'h00,8'h00}; // L
        Char_Matrix[13] = {8'h00,8'h00,8'h63,8'h77,8'h7F,8'h6B,8'h63,8'h63,8'h63,8'h63,8'h63,8'h63,8'h00,8'h00,8'h00,8'h00}; // M
        Char_Matrix[14] = {8'h00,8'h00,8'h63,8'h63,8'h73,8'h7B,8'h7F,8'h6F,8'h67,8'h63,8'h63,8'h63,8'h00,8'h00,8'h00,8'h00}; // N
        Char_Matrix[15] = {8'h00,8'h00,8'h1C,8'h36,8'h63,8'h63,8'h63,8'h63,8'h63,8'h63,8'h36,8'h1C,8'h00,8'h00,8'h00,8'h00}; // O
        Char_Matrix[16] = {8'h00,8'h00,8'h7E,8'h33,8'h33,8'h33,8'h3E,8'h30,8'h30,8'h30,8'h30,8'h78,8'h00,8'h00,8'h00,8'h00}; // P
        Char_Matrix[17] = {8'h00,8'h00,8'h3E,8'h63,8'h63,8'h63,8'h63,8'h63,8'h63,8'h6B,8'h6F,8'h3E,8'h06,8'h07,8'h00,8'h00}; // Q
        Char_Matrix[18] = {8'h00,8'h00,8'h7E,8'h33,8'h33,8'h33,8'h3E,8'h36,8'h36,8'h33,8'h33,8'h73,8'h00,8'h00,8'h00,8'h00}; // R
        Char_Matrix[19] = {8'h00,8'h00,8'h3E,8'h63,8'h63,8'h30,8'h1C,8'h06,8'h03,8'h63,8'h63,8'h3E,8'h00,8'h00,8'h00,8'h00}; // S
        Char_Matrix[20] = {8'h00,8'h00,8'hFF,8'hDB,8'h99,8'h18,8'h18,8'h18,8'h18,8'h18,8'h18,8'h3C,8'h00,8'h00,8'h00,8'h00}; // T
        Char_Matrix[21] = {8'h00,8'h00,8'h63,8'h63,8'h63,8'h63,8'h63,8'h63,8'h63,8'h63,8'h63,8'h3E,8'h00,8'h00,8'h00,8'h00}; // U
        Char_Matrix[22] = {8'h00,8'h00,8'h63,8'h63,8'h63,8'h63,8'h63,8'h63,8'h63,8'h36,8'h1C,8'h08,8'h00,8'h00,8'h00,8'h00}; // V
        Char_Matrix[23] = {8'h00,8'h00,8'h63,8'h63,8'h63,8'h63,8'h63,8'h6B,8'h6B,8'h7F,8'h36,8'h36,8'h00,8'h00,8'h00,8'h00}; // W
        Char_Matrix[24] = {8'h00,8'h00,8'hC3,8'hC3,8'h66,8'h3C,8'h18,8'h18,8'h3C,8'h66,8'hC3,8'hC3,8'h00,8'h00,8'h00,8'h00}; // X
        Char_Matrix[25] = {8'h00,8'h00,8'hC3,8'hC3,8'hC3,8'h66,8'h3C,8'h18,8'h18,8'h18,8'h18,8'h3C,8'h00,8'h00,8'h00,8'h00}; // Y
        Char_Matrix[26] = {8'h00,8'h00,8'h7F,8'h63,8'h43,8'h06,8'h0C,8'h18,8'h30,8'h61,8'h63,8'h7F,8'h00,8'h00,8'h00,8'h00}; // Z
        Char_Matrix[27] = {8'h00,8'h00,8'h00,8'h00,8'h00,8'h3C,8'h46,8'h06,8'h3E,8'h66,8'h66,8'h3B,8'h00,8'h00,8'h00,8'h00}; // a
        Char_Matrix[28] = {8'h00,8'h00,8'h70,8'h30,8'h30,8'h3C,8'h36,8'h33,8'h33,8'h33,8'h33,8'h6E,8'h00,8'h00,8'h00,8'h00}; // b
        Char_Matrix[29] = {8'h00,8'h00,8'h00,8'h00,8'h00,8'h3E,8'h63,8'h60,8'h60,8'h60,8'h63,8'h3E,8'h00,8'h00,8'h00,8'h00}; // c
        Char_Matrix[30] = {8'h00,8'h00,8'h0E,8'h06,8'h06,8'h1E,8'h36,8'h66,8'h66,8'h66,8'h66,8'h3B,8'h00,8'h00,8'h00,8'h00}; // d
        Char_Matrix[31] = {8'h00,8'h00,8'h00,8'h00,8'h00,8'h3E,8'h63,8'h63,8'h7E,8'h60,8'h63,8'h3E,8'h00,8'h00,8'h00,8'h00}; // e
        Char_Matrix[32] = {8'h00,8'h00,8'h1C,8'h36,8'h32,8'h30,8'h7C,8'h30,8'h30,8'h30,8'h30,8'h78,8'h00,8'h00,8'h00,8'h00}; // f
        Char_Matrix[33] = {8'h00,8'h00,8'h00,8'h00,8'h00,8'h3B,8'h66,8'h66,8'h66,8'h66,8'h3E,8'h06,8'h66,8'h3C,8'h00,8'h00}; // g
        Char_Matrix[34] = {8'h00,8'h00,8'h70,8'h30,8'h30,8'h36,8'h3B,8'h33,8'h33,8'h33,8'h33,8'h73,8'h00,8'h00,8'h00,8'h00}; // h
        Char_Matrix[35] = {8'h00,8'h00,8'h0C,8'h0C,8'h00,8'h1C,8'h0C,8'h0C,8'h0C,8'h0C,8'h0C,8'h1E,8'h00,8'h00,8'h00,8'h00}; // i
        Char_Matrix[36] = {8'h00,8'h00,8'h06,8'h06,8'h00,8'h0E,8'h06,8'h06,8'h06,8'h06,8'h06,8'h66,8'h66,8'h3C,8'h00,8'h00}; // j
        Char_Matrix[37] = {8'h00,8'h00,8'h70,8'h30,8'h30,8'h33,8'h33,8'h36,8'h3C,8'h36,8'h33,8'h73,8'h00,8'h00,8'h00,8'h00}; // k
        Char_Matrix[38] = {8'h00,8'h00,8'h1C,8'h0C,8'h0C,8'h0C,8'h0C,8'h0C,8'h0C,8'h0C,8'h0C,8'h1E,8'h00,8'h00,8'h00,8'h00}; // l
        Char_Matrix[39] = {8'h00,8'h00,8'h00,8'h00,8'h00,8'h6E,8'h7F,8'h6B,8'h6B,8'h6B,8'h6B,8'h6B,8'h00,8'h00,8'h00,8'h00}; // m
        Char_Matrix[40] = {8'h00,8'h00,8'h00,8'h00,8'h00,8'h6E,8'h33,8'h33,8'h33,8'h33,8'h33,8'h33,8'h00,8'h00,8'h00,8'h00}; // n
        Char_Matrix[41] = {8'h00,8'h00,8'h00,8'h00,8'h00,8'h3E,8'h63,8'h63,8'h63,8'h63,8'h63,8'h3E,8'h00,8'h00,8'h00,8'h00}; // o
        Char_Matrix[42] = {8'h00,8'h00,8'h00,8'h00,8'h00,8'h6E,8'h33,8'h33,8'h33,8'h33,8'h3E,8'h30,8'h30,8'h78,8'h00,8'h00}; // p
        Char_Matrix[43] = {8'h00,8'h00,8'h00,8'h00,8'h00,8'h3B,8'h66,8'h66,8'h66,8'h66,8'h3E,8'h06,8'h06,8'h0F,8'h00,8'h00}; // q
        Char_Matrix[44] = {8'h00,8'h00,8'h00,8'h00,8'h00,8'h6E,8'h3B,8'h33,8'h30,8'h30,8'h30,8'h78,8'h00,8'h00,8'h00,8'h00}; // r
        Char_Matrix[45] = {8'h00,8'h00,8'h00,8'h00,8'h00,8'h3E,8'h63,8'h38,8'h0E,8'h03,8'h63,8'h3E,8'h00,8'h00,8'h00,8'h00}; // s
        Char_Matrix[46] = {8'h00,8'h00,8'h08,8'h18,8'h18,8'h7E,8'h18,8'h18,8'h18,8'h18,8'h1B,8'h0E,8'h00,8'h00,8'h00,8'h00}; // t
        Char_Matrix[47] = {8'h00,8'h00,8'h00,8'h00,8'h00,8'h66,8'h66,8'h66,8'h66,8'h66,8'h66,8'h3B,8'h00,8'h00,8'h00,8'h00}; // u
        Char_Matrix[48] = {8'h00,8'h00,8'h00,8'h00,8'h00,8'h63,8'h63,8'h36,8'h36,8'h1C,8'h1C,8'h08,8'h00,8'h00,8'h00,8'h00}; // v
        Char_Matrix[49] = {8'h00,8'h00,8'h00,8'h00,8'h00,8'h63,8'h63,8'h63,8'h6B,8'h6B,8'h7F,8'h36,8'h00,8'h00,8'h00,8'h00}; // w
        Char_Matrix[50] = {8'h00,8'h00,8'h00,8'h00,8'h00,8'h63,8'h36,8'h1C,8'h1C,8'h1C,8'h36,8'h63,8'h00,8'h00,8'h00,8'h00}; // x
        Char_Matrix[51] = {8'h00,8'h00,8'h00,8'h00,8'h00,8'h63,8'h63,8'h63,8'h63,8'h63,8'h3F,8'h03,8'h06,8'h3C,8'h00,8'h00}; // y
        Char_Matrix[52] = {8'h00,8'h00,8'h00,8'h00,8'h00,8'h7F,8'h66,8'h0C,8'h18,8'h30,8'h63,8'h7F,8'h00,8'h00,8'h00,8'h00}; // z
        Char_Matrix[53] = {8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00}; // FO
    end
    
    wire [127:0] Matrix;
    assign Matrix = Char_Matrix[alph];
    always @(*)
    begin
        if((dcnt & 1) == 'b0)
            Point <= Matrix[127 - (8*dV + dH)]; //Char_Matrix���ǴӸ�λ����λ���
        else
            Point <= 'b0;
    end
endmodule
